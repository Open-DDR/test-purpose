//==============================================================================
// DDR2 Memory Controller
// 
// Description: Top-level DDR2 memory controller module
// Author: Open DDR Project
// Date: 2025
//==============================================================================

`include "ddr2_pkg.sv"

module ddr2_controller #(
    parameter DATA_WIDTH = 64,
    parameter ADDR_WIDTH = 32,
    parameter BANK_WIDTH = 3,
    parameter ROW_WIDTH  = 14,
    parameter COL_WIDTH  = 10
) (
    // Clock and Reset
    input  logic                    clk,
    input  logic                    rst_n,
    
    // AXI4 Interface
    input  logic [ADDR_WIDTH-1:0]  axi_awaddr,
    input  logic [7:0]              axi_awlen,
    input  logic [2:0]              axi_awsize,
    input  logic [1:0]              axi_awburst,
    input  logic                    axi_awvalid,
    output logic                    axi_awready,
    
    input  logic [DATA_WIDTH-1:0]  axi_wdata,
    input  logic [DATA_WIDTH/8-1:0] axi_wstrb,
    input  logic                    axi_wlast,
    input  logic                    axi_wvalid,
    output logic                    axi_wready,
    
    output logic [1:0]              axi_bresp,
    output logic                    axi_bvalid,
    input  logic                    axi_bready,
    
    input  logic [ADDR_WIDTH-1:0]  axi_araddr,
    input  logic [7:0]              axi_arlen,
    input  logic [2:0]              axi_arsize,
    input  logic [1:0]              axi_arburst,
    input  logic                    axi_arvalid,
    output logic                    axi_arready,
    
    output logic [DATA_WIDTH-1:0]  axi_rdata,
    output logic [1:0]              axi_rresp,
    output logic                    axi_rlast,
    output logic                    axi_rvalid,
    input  logic                    axi_rready,
    
    // DDR2 Physical Interface
    output logic                    ddr_ck_p,
    output logic                    ddr_ck_n,
    output logic                    ddr_cke,
    output logic                    ddr_cs_n,
    output logic                    ddr_ras_n,
    output logic                    ddr_cas_n,
    output logic                    ddr_we_n,
    output logic [BANK_WIDTH-1:0]  ddr_ba,
    output logic [ROW_WIDTH-1:0]   ddr_a,
    inout  wire  [DATA_WIDTH-1:0]  ddr_dq,
    inout  wire  [DATA_WIDTH/8-1:0] ddr_dqs_p,
    inout  wire  [DATA_WIDTH/8-1:0] ddr_dqs_n,
    output logic [DATA_WIDTH/8-1:0] ddr_dm,
    output logic                    ddr_odt
);

    import ddr2_pkg::*;

    // Internal signals
    logic [ADDR_WIDTH-1:0] decoded_addr;
    logic [BANK_WIDTH-1:0] bank_addr;
    logic [ROW_WIDTH-1:0]  row_addr;
    logic [COL_WIDTH-1:0]  col_addr;
    
    ctrl_state_t current_state, next_state;
    bank_state_t bank_states [2**BANK_WIDTH-1:0];
    
    // Command decoder
    ddr2_cmd_decoder u_cmd_decoder (
        .clk        (clk),
        .rst_n      (rst_n),
        .axi_addr   (axi_awvalid ? axi_awaddr : axi_araddr),
        .bank_addr  (bank_addr),
        .row_addr   (row_addr),
        .col_addr   (col_addr)
    );
    
    // Bank state machine
    ddr2_bank_fsm u_bank_fsm (
        .clk        (clk),
        .rst_n      (rst_n),
        .bank_addr  (bank_addr),
        .row_addr   (row_addr),
        .col_addr   (col_addr),
        .ddr_ras_n  (ddr_ras_n),
        .ddr_cas_n  (ddr_cas_n),
        .ddr_we_n   (ddr_we_n),
        .ddr_ba     (ddr_ba),
        .ddr_a      (ddr_a),
        .ddr_cs_n   (ddr_cs_n),
        .ddr_cke    (ddr_cke),
        .ddr_odt    (ddr_odt)
    );
    
    // PHY interface
    ddr2_phy u_phy (
        .clk        (clk),
        .rst_n      (rst_n),
        .ddr_ck_p   (ddr_ck_p),
        .ddr_ck_n   (ddr_ck_n),
        .ddr_dq     (ddr_dq),
        .ddr_dqs_p  (ddr_dqs_p),
        .ddr_dqs_n  (ddr_dqs_n),
        .ddr_dm     (ddr_dm)
    );
    
    // Refresh controller
    ddr2_refresh_ctrl u_refresh_ctrl (
        .clk        (clk),
        .rst_n      (rst_n),
        .refresh_req(/* refresh request logic */)
    );

endmodule
